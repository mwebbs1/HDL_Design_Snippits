module Four_Seven_Seg_Display(
    input clk,
    input [3:0]hex_1, hex_2, hex_3, hex_4,
    input dot_1, dot_2, dot_3, dot_4,
    output reg [3:0]an_out,
    output reg [6:0]seg_out,
    output dot_out
    );
    
    reg [1:0]select;
    wire pulse;
    wire [6:0]seg_1, seg_2, seg_3, seg_4;
    localparam FPS = 50; // Frames per second
    
    Clk_Divider_FPS #(.FPS(FPS*4)) clk2FPS(.clk(clk), .pulse(pulse));
    
    Seven_Segment_Display SSD1(.num(hex_1), .Display(seg_1));
    Seven_Segment_Display SSD2(.num(hex_2), .Display(seg_2));
    Seven_Segment_Display SSD3(.num(hex_3), .Display(seg_3));
    Seven_Segment_Display SSD4(.num(hex_4), .Display(seg_4));
    
    // Switch which number we are displaying 4 times per FPS
    always @(posedge clk)
        select <= (pulse == 1) ? select + 2'd1 : select;
    
    // output logic
    // switching order so that first number is on the left.
    always @(select)
        case(select)
            2'd0: begin seg_out <= seg_1; an_out <= 4'b1110; end
            2'd1: begin seg_out <= seg_2; an_out <= 4'b1101; end
            2'd2: begin seg_out <= seg_3; an_out <= 4'b1011; end
            2'd3: begin seg_out <= seg_4; an_out <= 4'b0111; end
        endcase
    
endmodule

module Seven_Segment_Display (
	input [3:0] num, 
	output reg [6:0] Display);
	
	// num is as binary number up to 15
	
	// Note: This implementation is for a common anode
	// 		Hence the ~
	always @(*)
		case (num)
			4'b0000: Display = ~7'b0111111; // 0
			4'b0001: Display = ~7'b0000110; // 1
			4'b0010: Display = ~7'b1011011; // 2
			4'b0011: Display = ~7'b1001111; // 3
			4'b0100: Display = ~7'b1100110; // 4
			4'b0101: Display = ~7'b1101101; // 5
			4'b0110: Display = ~7'b1111101; // 6
			4'b0111: Display = ~7'b0000111; // 7
			4'b1000: Display = ~7'b1111111; // 8
			4'b1001: Display = ~7'b1101111; // 9
			4'b1010: Display = ~7'b1110111; // A
			4'b1011: Display = ~7'b1111100; // b
			4'b1100: Display = ~7'b0111001; // C
			4'b1101: Display = ~7'b1011110; // d
			4'b1110: Display = ~7'b1111001; // E
			4'b1111: Display = ~7'b1110001; // F
			default: Display = ~7'b0000000; // 
		endcase
endmodule
